//************************* Copyright(c)2024, All rights reserved *********************
//                     __            Project name         : 
//                  \,`~"~` /        File name            : xxxxxxxx.v
//  .-=-.           /    . .\        Module name          : xxxxxxxx
// / .-. \          {  =    Y}=      Generated            : 2023-11-06 20:31:11
// _/   \ \          \      /        Last modified        : 2023-11-28 13:58:15
//       \ \        _/`'`'`b         Target Device        : XILINX 7A35T
//        \ `.__.-'`        \-._     Tool Versions        : Vivado 2022.1
//         |            '.__ `'-;_   Description          : 
//         |            _.' `'-.__)                         
//          \    ;_..--'/     //  \  
//          |   /  /   |     //    | Author               :    
//          \  \ \__)   \   //    /  E-Mail               : 
//           \__)        './/   .'   Company              : 
//                         `'-'`     Modification History :
//
// -----------------------------------------------------------------------------------
// |Have you noticed the cute kitten above？ She will bless you to write perfect code!|
// -----------------------------------------------------------------------------------
//
//*************************************************************************************

//*************************** Module, Parameters & Ports ******************************
module moduleName #(
    parameter P1 = 1,
              P2 = 2
) (
    input   [ W:0] I1,
    input   [ W:0] I2,
    output  [ W:0] O1,
    output  [ W:0] O2
);

//*************************** Module, Parameters & Ports ******************************
//*********************************** Localpatams *************************************
//************************************** Reg ******************************************
//************************************* Wire ******************************************
//************************************ Assign *****************************************
//************************************ Always *****************************************
//********************************** Instances ****************************************

endmodule

